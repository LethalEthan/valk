module main

fn main() {
	println('welcome to valk')
}