module packet.login

// clientbound packet 0x00
// pub struct CB_Disconnect {
// 	reason		Chat
// }